*Biblioteca de circuitos
*============inversor================================
.Subckt INV a out vdd gnd
	Mp1 vdd a out vdd PMOS l=16n w=64n 
	Mn1 out a gnd gnd NMOS l=16n w=32n 		
.Ends INV
*====================NAND==========================
.Subckt NAND a b out vdd gnd 
*rede pull up
	Mpa vdd a out vdd PMOS l=16n w=64n 
	Mpb vdd b out vdd PMOS l=16n w=64n 
*rede pull down
	Mna out a x gnd NMOS l=16n w=32n 
	Mnb x b gnd gnd NMOS l=16n w=32n 	
.Ends NAND

*======================NAND3===========================
.Subckt NAND3 a b c out vdd gnd
*rede pull up
	Mpa vdd a out vdd PMOS l=16n w=64n 
	Mpb vdd b out vdd PMOS l=16n w=64n 
	Mpc vdd c vdd vdd PMOS l=16n w=64n 

*rede pull down
	Mna out a x gnd NMOS l=16n w=32n 
	Mnb x b y gnd NMOS l=16n w=32n 
	Mnc y c gnd gnd NMOS l=16n w=32n 

.Ends NAND3
*====================NAND4============================
.Subckt NAND4 a b c d out vdd gnd
*rede pull up
	Mpa vdd a out vdd PMOS l=16n w=64n 
	Mpb vdd b out vdd PMOS l=16n w=64n 
	Mpc vdd c out vdd PMOS l=16n w=64n 
	Mpd vdd d out vdd PMOS l=16n w=64n 

*rede pull down
	Mna out a x gnd NMOS l=16n w=32n 
	Mnb x b y gnd NMOS l=16n w=32n 
	Mnc y c z gnd NMOS l=16n w=32n 
	Mnd z d gnd gnd NMOS l=16n w=32n 

.Ends NAND4
*====================NAND5============================
.Subckt NAND5 a b c d e out vdd gnd
*rede pull up
	Mpa vdd a out vdd PMOS l=16n w=64n 
	Mpb vdd b out vdd PMOS l=16n w=64n 
	Mpc vdd c out vdd PMOS l=16n w=64n 
	Mpd vdd d out vdd PMOS l=16n w=64n 
	Mpe vdd e out vdd PMOS l=16n w=64n 

*rede pull down
	Mna out a x gnd NMOS l=16n w=32n 
	Mnb x b y gnd NMOS l=16n w=32n 
	Mnc y c z gnd NMOS l=16n w=32n 
	Mnd z d z1 gnd NMOS l=16n w=32n 
	Mne z1 e gnd gnd NMOS l=16n w=32n 

.Ends NAND5
*===================AND==============================
.Subckt AND a b out vdd gnd 
	Xn2 a b s vdd gnd NAND
	Xinv s out vdd gnd INV
.Ends AND
*=====================AND3===============================
.Subckt AND3 a b c out vdd gnd
	Xn3 a b c s vdd gnd NAND3
	Xinv s out vdd gnd INV
.Ends AND3
*=============================AND4============================
.Subckt AND4 a b c d out vdd gnd
	Xn4 a b c d s vdd gnd NAND4
	Xinv s out vdd gnd INV
.Ends AND4
*=============================AND5============================
.Subckt AND5 a b c d e out vdd gnd
	Xn5 a b c d e s vdd gnd NAND5
	Xinv s out vdd gnd INV
.Ends AND5
*===================NOR2=================================
.Subckt NOR a b out vdd gnd
	Mp1 vdd a x vdd PMOS l=16n w=64n 
	Mp2 x b out vdd PMOS l=16n w=64n 

	Mn1 out a gnd gnd NMOS l=16n w=32n 
	Mn2 out b gnd gnd NMOS l=16n w=32n 
.Ends NOR
*======================NOR3=============================
.Subckt NOR3 a b c out vdd gnd
	Mp1 vdd a x vdd PMOS l=16n w=64n 
	Mp2 x b y vdd PMOS l=16n w=64n 
	Mp3 y c out vdd PMOS l=16n w=64n 


	Mn1 out a gnd gnd NMOS l=16n w=32n 
	Mn2 out b gnd gnd NMOS l=16n w=32n 
	Mn3 out c gnd gnd NMOS l=16n w=32n 
.Ends NOR3
*=======================NOR4===============================
.Subckt NOR4 a b c d out vdd gnd
	Mp1 vdd a x vdd PMOS l=16n w=64n 
	Mp2 x b y vdd PMOS l=16n w=64n 
	Mp3 y c z vdd PMOS l=16n w=64n 
	Mp4 z d out vdd PMOS l=16n w=64n 

	
	Mn1 out a gnd gnd NMOS l=16n w=32n 
	Mn2 out b gnd gnd NMOS l=16n w=32n 
	Mn3 out c gnd gnd NMOS l=16n w=32n 
	Mn4 out d gnd gnd NMOS l=16n w=32n 

.Ends NOR4
*=====================NOR5===============================
.Subckt NOR5 a b c d e out vdd gnd
	Mp1 vdd a x vdd PMOS l=16n w=64n 
	Mp2 x b y vdd PMOS l=16n w=64n 
	Mp3 y c z vdd PMOS l=16n w=64n 
	Mp4 z d m vdd PMOS l=16n w=64n 
	Mp5 m e out vdd PMOS l=16n w=64n 

	Mn1 out a gnd gnd NMOS l=16n w=32n 
	Mn2 out b gnd gnd NMOS l=16n w=32n 
	Mn3 out c gnd gnd NMOS l=16n w=32n 
	Mn4 out d gnd gnd NMOS l=16n w=32n 
	Mn5 out e gnd gnd NMOS l=16n w=32n 

.Ends NOR5
*=========================OR2============================
.Subckt OR a b out vdd gnd
	Xnor a b s vdd gnd NOR
	Xinv s out vdd gnd INV
.Ends OR

*==============================OR3=======================
.Subckt OR3 a b c out vdd gnd
	Xn3 a b c s vdd gnd NOR3
	Xi1 s out vdd gnd INV
.Ends OR3

*===============================OR4=======================
.Subckt OR4 a b c d out vdd gnd
	Xn4 a b c d s vdd gnd NOR4
	Xi1 s out vdd gnd INV
.Ends

*============================OR5============================
.Subckt OR5 a b c d e out vdd gnd
	Xn5 a b c d e s vdd gnd NOR5
	Xi1 s out vdd gnd INV
.Ends

*=================XOR====================================
.Subckt XOR a b out vdd gnd 
*instanciacao inversores
			Xinv1 a inva vdd gnd INV
			Xinv2 b invb vdd gnd INV
*====================REDE PULL UP=====================
*Esquerda=============================================
			Mp1 vdd invb nodo1 vdd PMOS L=16n W=64n 
			Mp2 nodo1 a out vdd PMOS L=16n W=64n 
*Direita=============================================
			Mp3 vdd b nodo2 vdd PMOS L=16n W=64n 
			Mp4 nodo2 inva out vdd PMOS L=16n W=64n 
*===============REDE PULL DOWN=======================
*Esquerda=============================================
			Mn1 out b nodo3 gnd NMOS L=16n W=32n 
			Mn2 nodo3 a gnd gnd NMOS L=16n W=32n 
*Direita=============================================
			Mn3 out invb nodo4 gnd NMOS L=16n W=32n 
			Mn4 nodo4 inva gnd gnd NMOS L=16n W=32n 								
.Ends XOR

*==============================HALF ADDER========================
.Subckt HA in1 in2 soma c vdd gnd
	Xxor in1 in2 soma vdd gnd XOR
	Xand in1 in2 c vdd gnd AND
.Ends HA

*=============Declaracao dos transistores do Somador CMOS=============
.param L = 16nm
.param Wp_FA= 64nm
.param Wn_FA =32nm

.subckt FA_CMOS cin a b soma cout vdd gnd
*---Pull-Up-----
Mp1 vdd a nodox1 vdd pmos L=L W=(2*Wp_FA)
Mp2 nodox1 b coutneg vdd pmos L=L W=(2*Wp_FA)

Mp3 vdd a nodox2 vdd pmos L=L W=(2*Wp_FA)
Mp4 vdd b nodox2 vdd pmos L=L W=(2*Wp_FA)
Mp5 nodox2 cin coutneg vdd pmos L=L W=(2*Wp_FA)

Mp6 vdd a nodox3 vdd pmos L=L W=(2*Wp_FA)
Mp7 vdd b nodox3 vdd pmos L=L W=(2*Wp_FA)
Mp8 vdd cin nodox3 vdd pmos L=L W=(2*Wp_FA)
Mp9 nodox3 coutneg somaneg vdd pmos L=L W=(2*Wp_FA)

Mp10 vdd a nodox4 vdd pmos L=L W=(3*Wp_FA)
Mp11 nodox4 b nodox5 vdd pmos L=L W=(3*Wp_FA)
Mp12 nodox5 cin somaneg vdd pmos L=L W=(3*Wp_FA)

Mp13 vdd somaneg soma vdd pmos L=L W=Wp_FA
Mp14 vdd coutneg cout vdd pmos L=L W=Wp_FA

*---Pull-Down-----
Mn1 nodox6 a gnd gnd nmos L=L W=(2*Wn_FA)
Mn2 coutneg b nodox6 gnd nmos L=L W=(2*Wn_FA)

Mn3 nodox7 a gnd gnd nmos L=L W=(2*Wn_FA)
Mn4 nodox7 b gnd gnd nmos L=L W=(2*Wn_FA)
Mn5 coutneg cin nodox7 gnd nmos L=L W=(2*Wn_FA)

Mn6 nodox8 a gnd gnd nmos L=L W=(2*Wn_FA)
Mn7 nodox8 b gnd gnd nmos L=L W=(2*Wn_FA)
Mn8 nodox8 cin gnd gnd nmos L=L W=(2*Wn_FA)
Mn9 somaneg coutneg nodox8 gnd nmos L=L W=(2*Wn_FA)

Mn10 nodox9 a gnd gnd nmos L=L W=(3*Wn_FA)
Mn11 nodox10 b nodox9 gnd nmos L=L W=(3*Wn_FA)
Mn12 somaneg cin nodox10 gnd nmos L=L W=(3*Wn_FA)

Mn13 soma somaneg gnd gnd nmos L=L W=Wn_FA
Mn14 cout coutneg gnd gnd nmos L=L W=Wn_FA
.ends FA_CMOS 
 
*=============================AXA2===========================
.subckt AXA2 cin a b soma cout vdd gnd
.param len = 16nm
.param wp = 64nm
.param wn = 32nm
    *Rede PMOS
        Mp1 vdd a co vdd PMOS w=wp l=len
        Mp2 vdd a sc1 vdd PMOS w=wp l=len
        Mp3 vdd b sc1 vdd PMOS w=wp l=len
        Mp4 sc1 co su vdd PMOS w=wp l=len
        Mp5 vdd cin su vdd PMOS w=wp l=len
    *Rede NMOS
        Mn1 co a gnd gnd NMOS w=wn l=len
        Mn2 su co sc2 gnd NMOS w=wn l=len
        Mn3 sc2 cin gnd gnd NMOS w=wn l=len
        Mn4 su cin sc3 gnd NMOS w=wn l=len
        Mn5 sc3 a sc4 gnd NMOS w=wn l=len
        Mn6 sc4 b gnd gnd NMOS w=wn l=len
Xcout co cout vdd gnd Inv
Xsum su soma vdd gnd Inv
.ends AXA2

*========CIRCUITO CAS======================================
.Subckt CAS cin yi sel enb pin soma cout vdd gnd
	Xxor sel yi a vdd gnd XOR
	Xand enb a b vdd gnd AND
	Xsum cin pin b soma cout vdd gnd FA_CMOS
.Ends CAS

*==========CAS AXA2====================================================
.Subckt CASAXA2 cin yi sel enb pin soma cout vdd gnd
	Xxor sel yi a vdd gnd XOR
	Xand enb a b vdd gnd AND
	Xsum cin pin b soma cout vdd gnd AXA2
.Ends CASAXA2


*====================WHITE CELL=================
.subckt whiteCell ci si a b soma cout vdd gnd
	Xand a b x vdd gnd AND
	Xsomador ci si x soma cout vdd gnd FA_CMOS
.ends whiteCell
 
*====================AXA2 WHITE CELL=================
.subckt WCAXA2 ci si a b soma cout vdd gnd
	Xand a b x vdd gnd AND
	Xsomador ci si x soma cout vdd gnd AXA2
.ends WCAXA2
 
 
*=====================GRAY CELL==============================
.subckt grayCell ci si a b soma cout vdd gnd
	Xnand a b x vdd gnd NAND
	Xsomador ci si x soma cout vdd gnd FA_CMOS
.ends grayCell
 
*=====================VEDIC 2===================================
.Subckt VEDIC2 ina0 ina1 inb0 inb1 p0 p1 p2 p3 vdd gnd
	Xand0 ina0 inb0 p0 vdd gnd AND
	Xand1 ina0 inb1 x0 vdd gnd AND 
	Xand2 ina1 inb0 x1 vdd gnd AND
	Xand3 ina1 inb1 x3 vdd gnd AND
	Xha1 x0 x1 p1 x2 vdd gnd HA
	Xha2 x2 x3 p2 p3 vdd gnd HA
.Ends VEDIC2 

*==============================CLA 4=================================
.Subckt CLA4 cin a0 a1 a2 a3 b0 b1 b2 b3 s0 s1 s2 s3 c4 PG GG vdd gnd
	Xx0 a0 b0 p0 vdd gnd OR
	Xx1 a1 b1 p1 vdd gnd OR
	Xx2 a2 b2 p2 vdd gnd OR
	Xx3 a3 b3 p3 vdd gnd OR
	Xa0 a0 b0 g0 vdd gnd AND
	Xa1 a1 b1 g1 vdd gnd AND
	Xa2 a2 b2 g2 vdd gnd AND
	Xa3 a3 b3 g3 vdd gnd AND
	
	Xand11 p0 cin nodo11 vdd gnd AND
	Xor1 g0 nodo11 c1 vdd gnd OR
	
	Xand21 g0 p1 nodo21 vdd gnd AND
	Xand22 cin p0 p1 nodo22 vdd gnd AND3
	Xor2 g1 nodo21 nodo22 c2 vdd gnd OR3
	
	Xand31 g1 p2 nodo31 vdd gnd AND
	Xand32 g0 p1 p2 nodo32 vdd gnd AND3
	Xand33 cin p0 p1 p2 nodo33 vdd gnd AND4
	Xor3 g2 nodo31 nodo32 nodo33 c3 vdd gnd OR4
	
	Xand41 g2 p3 nodo41 vdd gnd AND
	Xand42 g1 p2 p3 nodo42 vdd gnd AND3
	Xand43 g0 p1 p2 p3 nodo43 vdd gnd AND4
	Xand44 cin p0 p1 p2 p3 nodo44 vdd gnd AND5
	Xor4 g3 nodo41 nodo42 nodo43 nodo44 c4 vdd gnd OR5
	
	Xor_pg p0 p1 p2 p3 PG vdd gnd AND4
	Xor_gg g3 nodo41 nodo42 nodo43 GG vdd gnd OR4
		
	Xfa1 cin a0 b0 s0 cout1 vdd gnd FA_CMOS
	Xfa2 c1 a1 b1 s1 cout2 vdd gnd FA_CMOS
	Xfa3 c2 a2 b2 s2 cout3 vdd gnd FA_CMOS
	Xfa4 c3 a3 b3 s3 cout4 vdd gnd FA_CMOS
.Ends CLA4

*==============================RCA 4=================================
.Subckt RCA4 cin a0 a1 a2 a3 b0 b1 b2 b3 s0 s1 s2 s3 c4 vdd gnd
	Xfa1 cin a0 b0 s0 c1 vdd gnd FA_CMOS
	Xfa2 c1 a1 b1 s1 c2 vdd gnd FA_CMOS
	Xfa3 c2 a2 b2 s2 c3 vdd gnd FA_CMOS
	Xfa4 c3 a3 b3 s3 c4 vdd gnd FA_CMOS
.Ends RCA4

