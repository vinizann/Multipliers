*Biblioteca de circuitos
*============inversor================================
.Subckt INV a out vdd gnd
	Mp1 vdd a out vdd PMOS l=16n w=64n 
	Mn1 out a gnd gnd NMOS l=16n w=32n 		
.Ends INV
*====================NAND==========================
.Subckt NAND a b out vdd gnd 
*rede pull up
	Mpa vdd a out vdd PMOS l=16n w=64n 
	Mpb vdd b out vdd PMOS l=16n w=64n 
*rede pull down
	Mna out a x gnd NMOS l=16n w=32n 
	Mnb x b gnd gnd NMOS l=16n w=32n 	
.Ends NAND

*======================NAND3===========================
.Subckt NAND3 a b c out vdd gnd
*rede pull up
	Mpa vdd a out vdd PMOS l=16n w=64n 
	Mpb vdd b out vdd PMOS l=16n w=64n 
	Mpc vdd c vdd vdd PMOS l=16n w=64n 

*rede pull down
	Mna out a x gnd NMOS l=16n w=32n 
	Mnb x b y gnd NMOS l=16n w=32n 
	Mnc y c gnd gnd NMOS l=16n w=32n 

.Ends NAND3
*====================NAND4============================
.Subckt NAND4 a b c d out vdd gnd
*rede pull up
	Mpa vdd a out vdd PMOS l=16n w=64n 
	Mpb vdd b out vdd PMOS l=16n w=64n 
	Mpc vdd c out vdd PMOS l=16n w=64n 
	Mpd vdd d out vdd PMOS l=16n w=64n 

*rede pull down
	Mna out a x gnd NMOS l=16n w=32n 
	Mnb x b y gnd NMOS l=16n w=32n 
	Mnc y c z gnd NMOS l=16n w=32n 
	Mnd z d gnd gnd NMOS l=16n w=32n 

.Ends NAND4
*====================NAND5============================
.Subckt NAND5 a b c d e out vdd gnd
*rede pull up
	Mpa vdd a out vdd PMOS l=16n w=64n 
	Mpb vdd b out vdd PMOS l=16n w=64n 
	Mpc vdd c out vdd PMOS l=16n w=64n 
	Mpd vdd d out vdd PMOS l=16n w=64n 
	Mpe vdd e out vdd PMOS l=16n w=64n 

*rede pull down
	Mna out a x gnd NMOS l=16n w=32n 
	Mnb x b y gnd NMOS l=16n w=32n 
	Mnc y c z gnd NMOS l=16n w=32n 
	Mnd z d z1 gnd NMOS l=16n w=32n 
	Mne z1 e gnd gnd NMOS l=16n w=32n 

.Ends NAND5
*===================AND==============================
.Subckt AND a b out vdd gnd 
	Xn2 a b s vdd gnd NAND
	Xinv s out vdd gnd INV
.Ends AND
*=====================AND3===============================
.Subckt AND3 a b c out vdd gnd
	Xn3 a b c s vdd gnd NAND3
	Xinv s out vdd gnd INV
.Ends AND3
*=============================AND4============================
.Subckt AND4 a b c d out vdd gnd
	Xn4 a b c d s vdd gnd NAND4
	Xinv s out vdd gnd INV
.Ends AND4
*=============================AND5============================
.Subckt AND5 a b c d e out vdd gnd
	Xn5 a b c d e s vdd gnd NAND5
	Xinv s out vdd gnd INV
.Ends AND5
*===================NOR2=================================
.Subckt NOR a b out vdd gnd
	Mp1 vdd a x vdd PMOS l=16n w=64n 
	Mp2 x b out vdd PMOS l=16n w=64n 

	Mn1 out a gnd gnd NMOS l=16n w=32n 
	Mn2 out b gnd gnd NMOS l=16n w=32n 
.Ends NOR
*======================NOR3=============================
.Subckt NOR3 a b c out vdd gnd
	Mp1 vdd a x vdd PMOS l=16n w=64n 
	Mp2 x b y vdd PMOS l=16n w=64n 
	Mp3 y c out vdd PMOS l=16n w=64n 


	Mn1 out a gnd gnd NMOS l=16n w=32n 
	Mn2 out b gnd gnd NMOS l=16n w=32n 
	Mn3 out c gnd gnd NMOS l=16n w=32n 
.Ends NOR3
*=======================NOR4===============================
.Subckt NOR4 a b c d out vdd gnd
	Mp1 vdd a x vdd PMOS l=16n w=64n 
	Mp2 x b y vdd PMOS l=16n w=64n 
	Mp3 y c z vdd PMOS l=16n w=64n 
	Mp4 z d out vdd PMOS l=16n w=64n 

	
	Mn1 out a gnd gnd NMOS l=16n w=32n 
	Mn2 out b gnd gnd NMOS l=16n w=32n 
	Mn3 out c gnd gnd NMOS l=16n w=32n 
	Mn4 out d gnd gnd NMOS l=16n w=32n 

.Ends NOR4
*=====================NOR5===============================
.Subckt NOR5 a b c d e out vdd gnd
	Mp1 vdd a x vdd PMOS l=16n w=64n 
	Mp2 x b y vdd PMOS l=16n w=64n 
	Mp3 y c z vdd PMOS l=16n w=64n 
	Mp4 z d m vdd PMOS l=16n w=64n 
	Mp5 m e out vdd PMOS l=16n w=64n 

	Mn1 out a gnd gnd NMOS l=16n w=32n 
	Mn2 out b gnd gnd NMOS l=16n w=32n 
	Mn3 out c gnd gnd NMOS l=16n w=32n 
	Mn4 out d gnd gnd NMOS l=16n w=32n 
	Mn5 out e gnd gnd NMOS l=16n w=32n 

.Ends NOR5
*=========================OR2============================
.Subckt OR a b out vdd gnd
	Xnor a b s vdd gnd NOR
	Xinv s out vdd gnd INV
.Ends OR

*==============================OR3=======================
.Subckt OR3 a b c out vdd gnd
	Xn3 a b c s vdd gnd NOR3
	Xi1 s out vdd gnd INV
.Ends OR3

*===============================OR4=======================
.Subckt OR4 a b c d out vdd gnd
	Xn4 a b c d s vdd gnd NOR4
	Xi1 s out vdd gnd INV
.Ends

*============================OR5============================
.Subckt OR5 a b c d e out vdd gnd
	Xn5 a b c d e s vdd gnd NOR5
	Xi1 s out vdd gnd INV
.Ends

*=================XOR====================================
.Subckt XOR a b out vdd gnd 
*instanciacao inversores
			Xinv1 a inva vdd gnd INV
			Xinv2 b invb vdd gnd INV
*====================REDE PULL UP=====================
*Esquerda=============================================
			Mp1 vdd invb nodo1 vdd PMOS L=16n W=64n 
			Mp2 nodo1 a out vdd PMOS L=16n W=64n 
*Direita=============================================
			Mp3 vdd b nodo2 vdd PMOS L=16n W=64n 
			Mp4 nodo2 inva out vdd PMOS L=16n W=64n 
*===============REDE PULL DOWN=======================
*Esquerda=============================================
			Mn1 out b nodo3 gnd NMOS L=16n W=32n 
			Mn2 nodo3 a gnd gnd NMOS L=16n W=32n 
*Direita=============================================
			Mn3 out invb nodo4 gnd NMOS L=16n W=32n 
			Mn4 nodo4 inva gnd gnd NMOS L=16n W=32n 								
.Ends XOR

*==============================HALF ADDER========================
.Subckt HA in1 in2 soma c vdd gnd
	Xxor in1 in2 soma vdd gnd XOR
	Xand in1 in2 c vdd gnd AND
.Ends HA

*=============Declaracao dos transistores do Somador CMOS=============
.param L = 16nm
.param Wp_FA= 64nm
.param Wn_FA =32nm

.subckt FA_CMOS cin a b soma cout vdd gnd
*---Pull-Up-----
Mp1 vdd a nodox1 vdd pmos L=L W=(2*Wp_FA)
Mp2 nodox1 b coutneg vdd pmos L=L W=(2*Wp_FA)

Mp3 vdd a nodox2 vdd pmos L=L W=(2*Wp_FA)
Mp4 vdd b nodox2 vdd pmos L=L W=(2*Wp_FA)
Mp5 nodox2 cin coutneg vdd pmos L=L W=(2*Wp_FA)

Mp6 vdd a nodox3 vdd pmos L=L W=(2*Wp_FA)
Mp7 vdd b nodox3 vdd pmos L=L W=(2*Wp_FA)
Mp8 vdd cin nodox3 vdd pmos L=L W=(2*Wp_FA)
Mp9 nodox3 coutneg somaneg vdd pmos L=L W=(2*Wp_FA)

Mp10 vdd a nodox4 vdd pmos L=L W=(3*Wp_FA)
Mp11 nodox4 b nodox5 vdd pmos L=L W=(3*Wp_FA)
Mp12 nodox5 cin somaneg vdd pmos L=L W=(3*Wp_FA)

Mp13 vdd somaneg soma vdd pmos L=L W=Wp_FA
Mp14 vdd coutneg cout vdd pmos L=L W=Wp_FA

*---Pull-Down-----
Mn1 nodox6 a gnd gnd nmos L=L W=(2*Wn_FA)
Mn2 coutneg b nodox6 gnd nmos L=L W=(2*Wn_FA)

Mn3 nodox7 a gnd gnd nmos L=L W=(2*Wn_FA)
Mn4 nodox7 b gnd gnd nmos L=L W=(2*Wn_FA)
Mn5 coutneg cin nodox7 gnd nmos L=L W=(2*Wn_FA)

Mn6 nodox8 a gnd gnd nmos L=L W=(2*Wn_FA)
Mn7 nodox8 b gnd gnd nmos L=L W=(2*Wn_FA)
Mn8 nodox8 cin gnd gnd nmos L=L W=(2*Wn_FA)
Mn9 somaneg coutneg nodox8 gnd nmos L=L W=(2*Wn_FA)

Mn10 nodox9 a gnd gnd nmos L=L W=(3*Wn_FA)
Mn11 nodox10 b nodox9 gnd nmos L=L W=(3*Wn_FA)
Mn12 somaneg cin nodox10 gnd nmos L=L W=(3*Wn_FA)

Mn13 soma somaneg gnd gnd nmos L=L W=Wn_FA
Mn14 cout coutneg gnd gnd nmos L=L W=Wn_FA
.ends FA_CMOS 
 
*=============================COPY===========================
.Subckt COPY a b cin sum cout vdd gnd
	Xa a coutneg vdd gnd INV
	Xcoutneg coutneg cout vdd gnd INV
	Xb b sumneg vdd gnd INV
	Xsumneg sumneg sum vdd gnd INV
.ends COPY



